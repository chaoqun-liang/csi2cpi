
module csi2cpi_wrapper 
	#(
		parameter  NUM_RX_LANE = 2,
		parameter  RX_GEAR = 8,
		parameter  DATA_WIDTH = 48
	)
	(  
		// DPHY RX Submodule
		input  logic                        	clk_p_i,
		input  logic                        	clk_n_i,
		input  logic [NUM_RX_LANE - 1 : 0]	d_p_io,
		input  logic [NUM_RX_LANE - 1 : 0]	d_n_io,
		input  logic 						clk_byte_fr_i ,
		input  logic						reset_n_i ,
		input  logic 						reset_byte_n_i , 
		input  logic 						reset_byte_fr_n_i , 
		input  logic [5:0]					ref_dt_i ,     // reference data type . see tb
		input  logic 						tx_ready_i ,   // hmmmm can it be removed ? come back here dude
		input  logic 						pd_dphy_i ,    // only for hardened dphy block, i am going for hardened for now
		
		input  logic                         clk_pixel_i,
		input  logic                         pixel_rstn_i,
		output logic                         vsync_o ,
		output logic                         hsync_o ,
		output logic [DATA_WIDTH - 1:0]      pixel_o 
	);
		
			
		logic								axis_mtvalid ; 
		logic        [47:0]					axis_mtdata ; 
		logic								axis_stready ; 
		logic								axis_srstn;
		logic	 							clk_byte ;         // generated byte clock from dphy to latch internal parallel bate data from dphy_rx_wrap
		logic								clk_byte_hs ; 
        
		
		
		logic [NUM_RX_LANE -1 :0]           lp_d_rx_p ; 
		logic [NUM_RX_LANE - 1 :0]           lp_d_rx_n ; 
		logic [NUM_RX_LANE*RX_GEAR - 1 :0]   bd ;  // csi2(byte) data from parser
		
		
		logic 								sp_en ; // short packet enable
		logic 								lp_en ; // long packet enable 
		logic 								lp_av_en ; // a sad follower of lp_en, asserts when received long packets actually match the referred data type 
		logic 								hs_sync ; // successful detection of start sync code in data lanes
						
		
		myDphy rx_dphy(
			.axis_mtvalid_o		(axis_mtvalid ),
			.axis_mtdata_o		(axis_mtdata ),
			.axis_stready_i		(axis_stready ),
			.clk_byte_o			(clk_byte ),
			.clk_byte_hs_o		(clk_byte_hs ),
			.clk_byte_fr_i		(clk_byte_fr_i ),
			.reset_n_i			(reset_n_i ),
			.reset_byte_n_i  	(reset_byte_n_i ),
			.reset_byte_fr_n_i	(reset_byte_fr_n_i ),
			.clk_p_io			(clk_p_i ),
			.clk_n_io			(clk_n_i ),
			.d_p_io				(d_p_io ),
			.d_n_io				(d_n_io ),
			.lp_d_rx_p_o		(lp_d_rx_p ),
			.lp_d_rx_n_o		(lp_d_rx_n ),
			.bd_o				(bd ),
			.hs_sync_o			(hs_sync ),
			.ref_dt_i			(ref_dt_i ),
			.tx_rdy_i			(tx_ready_i ),
			.pd_dphy_i			(pd_dphy_i ),
			.sp_en_o			(sp_en ),
			.lp_en_o			(lp_en ),
			.lp_av_en_o			(lp_av_en )
			);
			

		axi4s_slave_if #(
			.DATA_WIDTH(DATA_WIDTH)
		) axi4s_slave ( 
			.axi4s_sclk_i       (clk_byte ),
			.axi4s_rstn_i       (axi4s_srstn ),
			.axi4s_svalid_i     (axis_mtvalid ),
			.axi4s_sready_o     (axis_stready ),
			.axi4s_sdata_i      (axis_mtdata)     // only take data type-5, word count-16 and payload-16. come back soon
			
		);
		
		
		sync_unpack sync_generator(
			.byte_clk_i			(clk_byte),
			.byte_rstn_i		(reset_n_i),
			.byte_vsync_i		(sp_en), // sp_en_o come back soon for a double check 
			.byte_hsync_i		(axis_mtvalid), // mtvalid_o shall work
			.pixel_clk_i		(clk_pixel_i),
			.pixel_rstn_i		(pixel_rstn_i),
			.vsync_o			(vsync_o),
			.hsync_o		    (hsync_o)						
	    );
	
	
		payload_unpack #(
			.DATA_WIDTH(DATA_WIDTH)
	   ) payload_generator (
			.byte_clk_i			(clk_byte),
			.byte_rstn_i		(reset_n_i),
			.pixel_clk_i		(clk_pixel_i),
			.pixel_rstn_i		(pixel_rstn_i),
			.wr_en_i			(),
			.rd_en_i			(),
			.vsync_o			(),
			.hsync_o			(),
			.wr_data_i			(),  // 16 LSB of trimmed mtdata 
			.rd_data_o			(pixel_o)					
     	);
	
	
endmodule			
		
